library verilog;
use verilog.vl_types.all;
entity multiMips is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end multiMips;
